module lstm_cell();//clk, rst, h_in, h_out);
//	parameter DATA_WIDTH = 16;
//	parameter FRACT_WIDTH = 8;
//	
//	input clk, rst;
//	
//	
//	// internal regs and wires
//	reg [DATA_WIDTH-1:0] C, h_prev;
//	
//	// f = sigmoid( WeightAndBias(  ) );
	
	
	
	
	
	


endmodule
